module add (a,b,c,sum);

input a,b,c;
output sum;

assign sum= a^b^c;

endmodule
