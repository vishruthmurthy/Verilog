`include "Register2.sv"
`include "Register1.sv"
`include "Adder.sv"
`include "Counter.sv"
`include "Comparator.sv"



